module hazard_detection_unit(
    input id_ex_memread,
    input [4:0] id_ex_rd,
    input [4:0] if_id_rs1,
    input [4:0] if_id_rs2,
    output pc_stall,
    output if_id_stall,
    output stall_mux
);







endmodule