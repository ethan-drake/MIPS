/CMC/kits/cadence/GPDK045/giolib045_v3.3/lef/giolib045.lef